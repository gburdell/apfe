module foo; i
/* block comment
with //line comment
*/
input foo; //line comment /*block comment*/
endmodule
