`define M 16
