`timescale  1ps/1ps
`ifndef N
`define N 4
`endif
`define N 5

module m1 (input [`N-1:0] d);
endmodule
