`define MM 12
