`include "m1.vh"

module m2;
endmodule
