`include "d.vh"

module m1;
endmodule
