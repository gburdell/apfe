`define PASTE /``/this is a comment
`PASTE
module m3;
`PASTE
endmodule
`undef DOOPY
`undef PASTE
