`define M 4