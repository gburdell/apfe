`line 1 "foo.v" 0
module g();
   a b(.c());
   a #1  b(.c());
endmodule
