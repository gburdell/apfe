module m2();
endmodule
