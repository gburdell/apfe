module m1(input p1, p2, output p3);
{ID1}; {ID2};
endmodule
